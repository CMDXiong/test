* 4 BIT ALU - 74LS181 EQUIV                     Revised:  December 29, 1996
* \ICED181\TOP181.SCH                           Revision: B
* P&D Engineering Consultants, Inc.
* 1970 Chalon Glen Court
* Livermore, CA  94550-8205
* Phone(510) 606-1285 /Fax (510) 606-1297
* 
.SUBCKT TOP181 VDD VSS A0 A1 A2 A3 B0 B1 B2 B3 S0 S1 S2 S3 M CN
+ GB CN4 PB F3B AEQB F2B F1B F0B
XINT1 VDD VSS M I INV3        
XINT3 VDD VSS 10059 AEQB INV3        
XNAT2 VDD VSS F3B F2B F1B F0B 10059 NAND4        
XXBIT3 A3 B3 A B S0 S1 S2 S3 VDD VSS ONEBIT
XXBIT2 A2 B2 C D S0 S1 S2 S3 VDD VSS ONEBIT
XXBIT1 A1 B1 E F S0 S1 S2 S3 VDD VSS ONEBIT
XXBIT0 A0 B0 G H S0 S1 S2 S3 VDD VSS ONEBIT
XXB0STF CN E F F0B F1B G H I VDD VSS B0STF
XXB1STF C CN D E F F2B G H I VDD VSS B1STF
XXB2STF A B C CN D E F F3B G H I VDD VSS B2STF
XXB3STF A B C CN CN4 D E F G GB H PB VDD VSS B3STF
.ENDS
.SUBCKT ONEBIT A B OT1 OT2 S0 S1 S2 S3 VDD VSS 
XIN1 VDD VSS B 10062 INV1        
XNA2 VDD VSS B S3 A 10055 NAND3        
XNA3 VDD VSS A S2 10062 10060 NAND3        
XNA4 VDD VSS 10055 10060 10058 NAND2        
XIN5 VDD VSS 10058 OT1 INV3        
XNA6 VDD VSS 10062 S1 10063 NAND2        
XNA7 VDD VSS S0 B 10065 NAND2        
XNA8 VDD VSS 10063 10065 A 10066 NAND3        
XIN9 VDD VSS 10066 OT2 INV3        
.ENDS
.SUBCKT B0STF CN E F F0B F1B G H I VDD VSS 
XXR0_1 VDD VSS E F 10071 XOR        
XXR0_2 VDD VSS 10071 10075 F1B XOR        
XNA0_3 VDD VSS CN G I 10078 NAND3        
XNA0_4 VDD VSS H I 10081 NAND2        
XNA0_5 VDD VSS 10078 10081 10080 NAND2        
XIN0_6 VDD VSS 10080 10075 INV1        
XXR0_7 VDD VSS H G 10083 XOR        
XXR0_8 VDD VSS 10083 10085 F0B XOR        
XNA0_9 VDD VSS CN I 10085 NAND2        
.ENDS
.SUBCKT B1STF C CN D E F F2B G H I VDD VSS 
XXR1_1 VDD VSS D C 10088 XOR        
XXR1_2 VDD VSS 10088 10092 F2B XOR        
XNA1_3 VDD VSS CN G E I 10095 NAND4        
XNA1_4 VDD VSS E H I 10099 NAND3        
XNA1_5 VDD VSS F I 10101 NAND2        
XNA1_6 VDD VSS 10095 10099 10101 10100 NAND3        
XIN1_7 VDD VSS 10100 10092 INV1        
.ENDS
.SUBCKT B2STF A B C CN D E F F3B G H I VDD VSS 
XXR2_1 VDD VSS B A 10108 XOR        
XNA2_3 VDD VSS CN G E C I 10116 NAND5        
XNA2_4 VDD VSS E C H I 10119 NAND4        
XNA2_5 VDD VSS C F I 10122 NAND3        
XNA2_6 VDD VSS D I 10123 NAND2        
XNA2_7 VDD VSS 10116 10119 10122 10123 10121 NAND4        
XIN2_8 VDD VSS 10121 10112 INV1        
XXR2_2 VDD VSS 10108 10112 F3B XOR        
.ENDS
.SUBCKT B3STF A B C CN CN4 D E F G GB H PB VDD VSS 
XIN3_1 VDD VSS B 10128 INV1        
XNA3_2 VDD VSS A D 10131 NAND2        
XNA3_3 VDD VSS A C F 10135 NAND3        
XNA3_4 VDD VSS A C E H 10136 NAND4        
XNA3_6 VDD VSS A C E G PB NAND4        
XNA3_8 VDD VSS 10128 10131 10135 10136 10133 NAND4        
XNA3_10 VDD VSS GB 10142 CN4 NAND2        
XIN3_9 VDD VSS 10133 GB INV3        
XNA3_5 VDD VSS A C E G CN 10142 NAND5        
.ENDS
.SUBCKT INV1 VDD VSS IN OUT 
MN1 OUT IN VSS VSS MN W=2U L=1.0U      
MP1 OUT IN VDD VDD MP W=4U L=1.0U      
.ENDS
.SUBCKT INV3 VDD VSS IN OUT
MN1 OUT IN VSS VSS MN W=6U L=1.0U      
MP1 OUT IN VDD VDD MP W=12U L=1.0U      
.ENDS
.SUBCKT NAND2 VDD VSS IN1 IN2 OUT 
MP2 OUT IN2 VDD VDD MP W=4U L=1.0U      
MP1 OUT IN1 VDD VDD MP W=4U L=1.0U      
MN1 OUT IN1 10091 VSS MN W=2U L=1.0U      
MN2 10091 IN2 VSS VSS MN W=2U L=1.0U      
.ENDS
.SUBCKT NAND3 VDD VSS IN1 IN2 IN3 OUT 
MP3 OUT IN3 VDD VDD MP W=4U L=1.0U      
MP2 OUT IN2 VDD VDD MP W=4U L=1.0U      
MP1 OUT IN1 VDD VDD MP W=4U L=1.0U      
MN1 OUT IN1 10086 VSS MN W=3U L=1.0U      
MN2 10086 IN2 10087 VSS MN W=3U L=1.0U      
MN3 10087 IN3 VSS VSS MN W=3U L=1.0U      
.ENDS
.SUBCKT NAND4 VDD VSS IN1 IN2 IN3 IN4 OUT 
MN4 10113 IN4 VSS VSS MN W=4.0U L=1.0U      
MN3 10112 IN3 10113 VSS MN W=4.0U L=1.0U      
MN2 10111 IN2 10112 VSS MN W=4.0U L=1.0U      
MN1 OUT IN1 10111 VSS MN W=4.0U L=1.0U      
MP1 OUT IN1 VDD VDD MP W=4.0U L=1.0U      
MP2 OUT IN2 VDD VDD MP W=4.0U L=1.0U      
MP3 OUT IN3 VDD VDD MP W=4.0U L=1.0U      
MP4 OUT IN4 VDD VDD MP W=4.0U L=1.0U      
.ENDS
.SUBCKT NAND5 VDD VSS IN1 IN2 IN3 IN4 IN5 OUT 
MN4 10244 IN4 10245 VSS MN W=4.0U L=1.0U      
MN3 10243 IN3 10244 VSS MN W=4.0U L=1.0U      
MN2 10242 IN2 10243 VSS MN W=4.0U L=1.0U      
MN1 OUT IN1 10242 VSS MN W=4.0U L=1.0U      
MP1 OUT IN1 VDD VDD MP W=4.0U L=1.0U      
MP2 OUT IN2 VDD VDD MP W=4.0U L=1.0U      
MP3 OUT IN3 VDD VDD MP W=4.0U L=1.0U      
MP4 OUT IN4 VDD VDD MP W=4.0U L=1.0U      
MN5 10245 IN5 VSS VSS MN W=4.0U L=1.0U      
MP5 OUT IN5 VDD VDD MP W=4.0U L=1.0U      
.ENDS
.SUBCKT XOR VDD VSS IN1 IN2 OUT 
MN1 10148 IN1 VSS VSS MN W=3U L=1.0U      
MN2 10152 10148 VSS VSS MN W=2U L=1.0U      
MN4 OUT IN2 10148 VSS MN W=2U L=1.0U      
MN5 OUT 10149 10152 VSS MN W=4U L=1.0U      
MN3 10149 IN2 VSS VSS MN W=2U L=1.0U      
MP2 10149 IN2 VDD VDD MP W=4U L=1.0U      
MP1 10148 IN1 VDD VDD MP W=5U L=1.0U      
MP3 OUT 10149 10148 VDD MP W=5U L=1.0U      
MP4 OUT 10148 10149 VDD MP W=6U L=1.0U      
.ENDS
.END
